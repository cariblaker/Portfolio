module state_machine(

);


endmodule 