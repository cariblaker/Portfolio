module myBCDAdder(
	input [3:0]a,
	input [3:0]b,
	output [7:0]X
);


	assign X = ( (a + b) < 10 ) ? (a + b) : ( (a + b) == 10 ) ? 8'b00010000 : ( (a + b) == 11 ) ? 8'b00010001 : ((a + b) == 12) ? 8'b00010010 : ((a + b) == 13) ? 8'b00010011 : ((a + b) == 14) ? 8'b00010100 : ((a + b) == 15) ? 8'b00010101 : ((a + b) == 16) ? 8'b00010110 : ((a + b) == 17) ? 8'b00010111 : 8'b00011000;

endmodule
