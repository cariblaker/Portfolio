module row(
	input clk,
	output reg [3:0]rout
);





endmodule 
