module my_modu(
	input sx,
	input a,
	input b,
	output m_out
);


//wire [2:1]G;

//and U1(sx, G[1], G[2]);


endmodule